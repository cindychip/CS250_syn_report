VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram8t17x64
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 55.264 BY 52.288 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
  END O1[28]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
  END O1[32]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
  END O1[36]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
  END O1[40]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
  END O1[44]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
  END O1[48]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
  END O1[52]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
  END O1[56]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
  END O1[60]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.112 45.752 55.264 45.904 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.112 45.752 55.264 45.904 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.112 45.752 55.264 45.904 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.112 45.752 55.264 45.904 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.112 42.104 55.264 42.256 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.112 42.104 55.264 42.256 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.112 42.104 55.264 42.256 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.112 42.104 55.264 42.256 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.112 38.456 55.264 38.608 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.112 38.456 55.264 38.608 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.112 38.456 55.264 38.608 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.112 38.456 55.264 38.608 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.112 34.808 55.264 34.960 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.112 34.808 55.264 34.960 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.112 34.808 55.264 34.960 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.112 34.808 55.264 34.960 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.112 31.160 55.264 31.312 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.112 31.160 55.264 31.312 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.112 31.160 55.264 31.312 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.112 31.160 55.264 31.312 ;
    END
  END A1[4]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.584 0.000 3.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.584 0.000 3.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.584 0.000 3.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.584 0.000 3.736 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.888 0.000 4.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 3.888 0.000 4.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.888 0.000 4.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 3.888 0.000 4.040 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.192 0.000 4.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.192 0.000 4.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.192 0.000 4.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.192 0.000 4.344 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.496 0.000 4.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.496 0.000 4.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.496 0.000 4.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.496 0.000 4.648 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.800 0.000 4.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.800 0.000 4.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.800 0.000 4.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.800 0.000 4.952 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.104 0.000 5.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.104 0.000 5.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.104 0.000 5.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.104 0.000 5.256 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.408 0.000 5.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.408 0.000 5.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.408 0.000 5.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.408 0.000 5.560 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 5.712 0.000 5.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.712 0.000 5.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 5.712 0.000 5.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.712 0.000 5.864 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.016 0.000 6.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.016 0.000 6.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.016 0.000 6.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.016 0.000 6.168 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.320 0.000 6.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.320 0.000 6.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.320 0.000 6.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.320 0.000 6.472 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.624 0.000 6.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.624 0.000 6.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.624 0.000 6.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.624 0.000 6.776 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.928 0.000 7.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.928 0.000 7.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.928 0.000 7.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.928 0.000 7.080 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.232 0.000 7.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.232 0.000 7.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.232 0.000 7.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.232 0.000 7.384 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.536 0.000 7.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.536 0.000 7.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.536 0.000 7.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.536 0.000 7.688 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.840 0.000 7.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.840 0.000 7.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.840 0.000 7.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.840 0.000 7.992 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.144 0.000 8.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.144 0.000 8.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.144 0.000 8.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.144 0.000 8.296 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.448 0.000 8.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.448 0.000 8.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.448 0.000 8.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.448 0.000 8.600 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.752 0.000 8.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.752 0.000 8.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.752 0.000 8.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.752 0.000 8.904 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.056 0.000 9.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.056 0.000 9.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.056 0.000 9.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.056 0.000 9.208 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.360 0.000 9.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.360 0.000 9.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.360 0.000 9.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.360 0.000 9.512 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.664 0.000 9.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.664 0.000 9.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.664 0.000 9.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.664 0.000 9.816 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.968 0.000 10.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.968 0.000 10.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.968 0.000 10.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.968 0.000 10.120 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.272 0.000 10.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.272 0.000 10.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.272 0.000 10.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.272 0.000 10.424 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.576 0.000 10.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.576 0.000 10.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.576 0.000 10.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.576 0.000 10.728 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.880 0.000 11.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.880 0.000 11.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.880 0.000 11.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.880 0.000 11.032 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.184 0.000 11.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.184 0.000 11.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.184 0.000 11.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.184 0.000 11.336 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.488 0.000 11.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.488 0.000 11.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.488 0.000 11.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.488 0.000 11.640 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.792 0.000 11.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.792 0.000 11.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.792 0.000 11.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.792 0.000 11.944 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.096 0.000 12.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.096 0.000 12.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.096 0.000 12.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.096 0.000 12.248 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.400 0.000 12.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.400 0.000 12.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.400 0.000 12.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.400 0.000 12.552 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.704 0.000 12.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.704 0.000 12.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.704 0.000 12.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.704 0.000 12.856 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.008 0.000 13.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.008 0.000 13.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.008 0.000 13.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.008 0.000 13.160 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.312 0.000 13.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.312 0.000 13.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.312 0.000 13.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.312 0.000 13.464 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.616 0.000 13.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.616 0.000 13.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.616 0.000 13.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.616 0.000 13.768 0.152 ;
    END
  END I2[31]

  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.920 0.000 14.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.920 0.000 14.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.920 0.000 14.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.920 0.000 14.072 0.152 ;
    END
  END I2[32]

  PIN I2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.224 0.000 14.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.224 0.000 14.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.224 0.000 14.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.224 0.000 14.376 0.152 ;
    END
  END I2[33]

  PIN I2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.528 0.000 14.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.528 0.000 14.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.528 0.000 14.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.528 0.000 14.680 0.152 ;
    END
  END I2[34]

  PIN I2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.832 0.000 14.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.832 0.000 14.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.832 0.000 14.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.832 0.000 14.984 0.152 ;
    END
  END I2[35]

  PIN I2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.136 0.000 15.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.136 0.000 15.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.136 0.000 15.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.136 0.000 15.288 0.152 ;
    END
  END I2[36]

  PIN I2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.440 0.000 15.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.440 0.000 15.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.440 0.000 15.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.440 0.000 15.592 0.152 ;
    END
  END I2[37]

  PIN I2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.744 0.000 15.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.744 0.000 15.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.744 0.000 15.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.744 0.000 15.896 0.152 ;
    END
  END I2[38]

  PIN I2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.048 0.000 16.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.048 0.000 16.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.048 0.000 16.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.048 0.000 16.200 0.152 ;
    END
  END I2[39]

  PIN I2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.352 0.000 16.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.352 0.000 16.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.352 0.000 16.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.352 0.000 16.504 0.152 ;
    END
  END I2[40]

  PIN I2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.656 0.000 16.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.656 0.000 16.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.656 0.000 16.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.656 0.000 16.808 0.152 ;
    END
  END I2[41]

  PIN I2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.960 0.000 17.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.960 0.000 17.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.960 0.000 17.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.960 0.000 17.112 0.152 ;
    END
  END I2[42]

  PIN I2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.264 0.000 17.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.264 0.000 17.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.264 0.000 17.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.264 0.000 17.416 0.152 ;
    END
  END I2[43]

  PIN I2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.568 0.000 17.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.568 0.000 17.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.568 0.000 17.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.568 0.000 17.720 0.152 ;
    END
  END I2[44]

  PIN I2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.872 0.000 18.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.872 0.000 18.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.872 0.000 18.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.872 0.000 18.024 0.152 ;
    END
  END I2[45]

  PIN I2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.176 0.000 18.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.176 0.000 18.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.176 0.000 18.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.176 0.000 18.328 0.152 ;
    END
  END I2[46]

  PIN I2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.480 0.000 18.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.480 0.000 18.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.480 0.000 18.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.480 0.000 18.632 0.152 ;
    END
  END I2[47]

  PIN I2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.784 0.000 18.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.784 0.000 18.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.784 0.000 18.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.784 0.000 18.936 0.152 ;
    END
  END I2[48]

  PIN I2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.088 0.000 19.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.088 0.000 19.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.088 0.000 19.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.088 0.000 19.240 0.152 ;
    END
  END I2[49]

  PIN I2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.392 0.000 19.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.392 0.000 19.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.392 0.000 19.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.392 0.000 19.544 0.152 ;
    END
  END I2[50]

  PIN I2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.696 0.000 19.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.696 0.000 19.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.696 0.000 19.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.696 0.000 19.848 0.152 ;
    END
  END I2[51]

  PIN I2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.000 0.000 20.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.000 0.000 20.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.000 0.000 20.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.000 0.000 20.152 0.152 ;
    END
  END I2[52]

  PIN I2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.304 0.000 20.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.304 0.000 20.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.304 0.000 20.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.304 0.000 20.456 0.152 ;
    END
  END I2[53]

  PIN I2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.608 0.000 20.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.608 0.000 20.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.608 0.000 20.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.608 0.000 20.760 0.152 ;
    END
  END I2[54]

  PIN I2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.912 0.000 21.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.912 0.000 21.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.912 0.000 21.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.912 0.000 21.064 0.152 ;
    END
  END I2[55]

  PIN I2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.216 0.000 21.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.216 0.000 21.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.216 0.000 21.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.216 0.000 21.368 0.152 ;
    END
  END I2[56]

  PIN I2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.520 0.000 21.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.520 0.000 21.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.520 0.000 21.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.520 0.000 21.672 0.152 ;
    END
  END I2[57]

  PIN I2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.824 0.000 21.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.824 0.000 21.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.824 0.000 21.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.824 0.000 21.976 0.152 ;
    END
  END I2[58]

  PIN I2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.128 0.000 22.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.128 0.000 22.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.128 0.000 22.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.128 0.000 22.280 0.152 ;
    END
  END I2[59]

  PIN I2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.432 0.000 22.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.432 0.000 22.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.432 0.000 22.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.432 0.000 22.584 0.152 ;
    END
  END I2[60]

  PIN I2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.736 0.000 22.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.736 0.000 22.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.736 0.000 22.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.736 0.000 22.888 0.152 ;
    END
  END I2[61]

  PIN I2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.040 0.000 23.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.040 0.000 23.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.040 0.000 23.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.040 0.000 23.192 0.152 ;
    END
  END I2[62]

  PIN I2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.344 0.000 23.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.344 0.000 23.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.344 0.000 23.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.344 0.000 23.496 0.152 ;
    END
  END I2[63]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 45.752 0.152 45.904 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 45.752 0.152 45.904 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 45.752 0.152 45.904 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 45.752 0.152 45.904 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 42.104 0.152 42.256 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 42.104 0.152 42.256 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 42.104 0.152 42.256 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 42.104 0.152 42.256 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 38.456 0.152 38.608 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 38.456 0.152 38.608 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 38.456 0.152 38.608 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 38.456 0.152 38.608 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 34.808 0.152 34.960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 34.808 0.152 34.960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 34.808 0.152 34.960 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 34.808 0.152 34.960 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 31.160 0.152 31.312 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 31.160 0.152 31.312 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 31.160 0.152 31.312 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 31.160 0.152 31.312 ;
    END
  END A2[4]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 13.072 0.152 13.224 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 13.072 0.152 13.224 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 13.072 0.152 13.224 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 13.072 0.152 13.224 ;
    END
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 50.288 7.195 52.288 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 50.288 7.195 52.288 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 50.288 7.195 52.288 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 50.288 9.915 52.288 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 50.288 9.915 52.288 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 50.288 9.915 52.288 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 51.984 0.000 55.264 0.304 ;
      RECT 51.680 0.000 51.528 0.304 ;
      RECT 51.376 0.000 51.224 0.304 ;
      RECT 51.072 0.000 50.920 0.304 ;
      RECT 49.856 0.000 49.704 0.304 ;
      RECT 48.640 0.000 48.488 0.304 ;
      RECT 47.424 0.000 47.272 0.304 ;
      RECT 46.208 0.000 46.056 0.304 ;
      RECT 44.992 0.000 44.840 0.304 ;
      RECT 43.776 0.000 43.624 0.304 ;
      RECT 42.560 0.000 42.408 0.304 ;
      RECT 41.344 0.000 41.192 0.304 ;
      RECT 40.128 0.000 39.976 0.304 ;
      RECT 38.912 0.000 38.760 0.304 ;
      RECT 37.696 0.000 37.544 0.304 ;
      RECT 36.480 0.000 36.328 0.304 ;
      RECT 35.264 0.000 35.112 0.304 ;
      RECT 34.048 0.000 33.896 0.304 ;
      RECT 32.832 0.000 32.680 0.304 ;
      RECT 54.960 46.056 55.264 50.136 ;
      RECT 54.960 42.408 55.264 45.600 ;
      RECT 54.960 38.760 55.264 41.952 ;
      RECT 54.960 35.112 55.264 38.304 ;
      RECT 54.960 31.464 55.264 34.656 ;
      RECT 54.960 13.376 55.264 31.008 ;
      RECT 54.960 0.304 55.264 12.920 ;
      RECT 0.000 0.000 3.432 0.304 ;
      RECT 3.888 0.000 3.736 0.304 ;
      RECT 4.192 0.000 4.040 0.304 ;
      RECT 5.408 0.000 5.256 0.304 ;
      RECT 6.624 0.000 6.472 0.304 ;
      RECT 7.840 0.000 7.688 0.304 ;
      RECT 9.056 0.000 8.904 0.304 ;
      RECT 10.272 0.000 10.120 0.304 ;
      RECT 11.488 0.000 11.336 0.304 ;
      RECT 12.704 0.000 12.552 0.304 ;
      RECT 13.920 0.000 13.768 0.304 ;
      RECT 15.136 0.000 14.984 0.304 ;
      RECT 16.352 0.000 16.200 0.304 ;
      RECT 17.568 0.000 17.416 0.304 ;
      RECT 18.784 0.000 18.632 0.304 ;
      RECT 20.000 0.000 19.848 0.304 ;
      RECT 21.216 0.000 21.064 0.304 ;
      RECT 22.432 0.000 22.280 0.304 ;
      RECT 23.648 0.000 31.464 0.304 ;
      RECT 0.000 46.056 0.304 50.136 ;
      RECT 0.000 42.408 0.304 45.600 ;
      RECT 0.000 38.760 0.304 41.952 ;
      RECT 0.000 35.112 0.304 38.304 ;
      RECT 0.000 31.464 0.304 34.656 ;
      RECT 0.000 13.376 0.304 31.008 ;
      RECT 0.000 0.304 0.304 12.920 ;
      RECT 0.000 50.136 5.043 52.288 ;
      RECT 7.355 50.136 7.763 52.288 ;
      RECT 10.067 50.136 55.264 52.288 ;
      RECT 0.304 0.304 54.960 50.136 ;
    LAYER M3 ;
      RECT 51.984 0.000 55.264 0.304 ;
      RECT 51.680 0.000 51.528 0.304 ;
      RECT 51.376 0.000 51.224 0.304 ;
      RECT 51.072 0.000 50.920 0.304 ;
      RECT 49.856 0.000 49.704 0.304 ;
      RECT 48.640 0.000 48.488 0.304 ;
      RECT 47.424 0.000 47.272 0.304 ;
      RECT 46.208 0.000 46.056 0.304 ;
      RECT 44.992 0.000 44.840 0.304 ;
      RECT 43.776 0.000 43.624 0.304 ;
      RECT 42.560 0.000 42.408 0.304 ;
      RECT 41.344 0.000 41.192 0.304 ;
      RECT 40.128 0.000 39.976 0.304 ;
      RECT 38.912 0.000 38.760 0.304 ;
      RECT 37.696 0.000 37.544 0.304 ;
      RECT 36.480 0.000 36.328 0.304 ;
      RECT 35.264 0.000 35.112 0.304 ;
      RECT 34.048 0.000 33.896 0.304 ;
      RECT 32.832 0.000 32.680 0.304 ;
      RECT 54.960 46.056 55.264 50.136 ;
      RECT 54.960 42.408 55.264 45.600 ;
      RECT 54.960 38.760 55.264 41.952 ;
      RECT 54.960 35.112 55.264 38.304 ;
      RECT 54.960 31.464 55.264 34.656 ;
      RECT 54.960 13.376 55.264 31.008 ;
      RECT 54.960 0.304 55.264 12.920 ;
      RECT 0.000 0.000 3.432 0.304 ;
      RECT 3.888 0.000 3.736 0.304 ;
      RECT 4.192 0.000 4.040 0.304 ;
      RECT 5.408 0.000 5.256 0.304 ;
      RECT 6.624 0.000 6.472 0.304 ;
      RECT 7.840 0.000 7.688 0.304 ;
      RECT 9.056 0.000 8.904 0.304 ;
      RECT 10.272 0.000 10.120 0.304 ;
      RECT 11.488 0.000 11.336 0.304 ;
      RECT 12.704 0.000 12.552 0.304 ;
      RECT 13.920 0.000 13.768 0.304 ;
      RECT 15.136 0.000 14.984 0.304 ;
      RECT 16.352 0.000 16.200 0.304 ;
      RECT 17.568 0.000 17.416 0.304 ;
      RECT 18.784 0.000 18.632 0.304 ;
      RECT 20.000 0.000 19.848 0.304 ;
      RECT 21.216 0.000 21.064 0.304 ;
      RECT 22.432 0.000 22.280 0.304 ;
      RECT 23.648 0.000 31.464 0.304 ;
      RECT 0.000 46.056 0.304 50.136 ;
      RECT 0.000 42.408 0.304 45.600 ;
      RECT 0.000 38.760 0.304 41.952 ;
      RECT 0.000 35.112 0.304 38.304 ;
      RECT 0.000 31.464 0.304 34.656 ;
      RECT 0.000 13.376 0.304 31.008 ;
      RECT 0.000 0.304 0.304 12.920 ;
      RECT 0.000 50.136 5.043 52.288 ;
      RECT 7.355 50.136 7.763 52.288 ;
      RECT 10.067 50.136 55.264 52.288 ;
      RECT 0.304 0.304 54.960 50.136 ;
    LAYER M4 ;
      RECT 51.984 0.000 55.264 0.304 ;
      RECT 51.680 0.000 51.528 0.304 ;
      RECT 51.376 0.000 51.224 0.304 ;
      RECT 51.072 0.000 50.920 0.304 ;
      RECT 49.856 0.000 49.704 0.304 ;
      RECT 48.640 0.000 48.488 0.304 ;
      RECT 47.424 0.000 47.272 0.304 ;
      RECT 46.208 0.000 46.056 0.304 ;
      RECT 44.992 0.000 44.840 0.304 ;
      RECT 43.776 0.000 43.624 0.304 ;
      RECT 42.560 0.000 42.408 0.304 ;
      RECT 41.344 0.000 41.192 0.304 ;
      RECT 40.128 0.000 39.976 0.304 ;
      RECT 38.912 0.000 38.760 0.304 ;
      RECT 37.696 0.000 37.544 0.304 ;
      RECT 36.480 0.000 36.328 0.304 ;
      RECT 35.264 0.000 35.112 0.304 ;
      RECT 34.048 0.000 33.896 0.304 ;
      RECT 32.832 0.000 32.680 0.304 ;
      RECT 54.960 46.056 55.264 50.136 ;
      RECT 54.960 42.408 55.264 45.600 ;
      RECT 54.960 38.760 55.264 41.952 ;
      RECT 54.960 35.112 55.264 38.304 ;
      RECT 54.960 31.464 55.264 34.656 ;
      RECT 54.960 13.376 55.264 31.008 ;
      RECT 54.960 0.304 55.264 12.920 ;
      RECT 0.000 0.000 3.432 0.304 ;
      RECT 3.888 0.000 3.736 0.304 ;
      RECT 4.192 0.000 4.040 0.304 ;
      RECT 5.408 0.000 5.256 0.304 ;
      RECT 6.624 0.000 6.472 0.304 ;
      RECT 7.840 0.000 7.688 0.304 ;
      RECT 9.056 0.000 8.904 0.304 ;
      RECT 10.272 0.000 10.120 0.304 ;
      RECT 11.488 0.000 11.336 0.304 ;
      RECT 12.704 0.000 12.552 0.304 ;
      RECT 13.920 0.000 13.768 0.304 ;
      RECT 15.136 0.000 14.984 0.304 ;
      RECT 16.352 0.000 16.200 0.304 ;
      RECT 17.568 0.000 17.416 0.304 ;
      RECT 18.784 0.000 18.632 0.304 ;
      RECT 20.000 0.000 19.848 0.304 ;
      RECT 21.216 0.000 21.064 0.304 ;
      RECT 22.432 0.000 22.280 0.304 ;
      RECT 23.648 0.000 31.464 0.304 ;
      RECT 0.000 46.056 0.304 50.136 ;
      RECT 0.000 42.408 0.304 45.600 ;
      RECT 0.000 38.760 0.304 41.952 ;
      RECT 0.000 35.112 0.304 38.304 ;
      RECT 0.000 31.464 0.304 34.656 ;
      RECT 0.000 13.376 0.304 31.008 ;
      RECT 0.000 0.304 0.304 12.920 ;
      RECT 0.000 50.136 5.043 52.288 ;
      RECT 7.355 50.136 7.763 52.288 ;
      RECT 10.067 50.136 55.264 52.288 ;
      RECT 0.304 0.304 54.960 50.136 ;
    LAYER M5 ;
      RECT 51.984 0.000 55.264 0.304 ;
      RECT 51.680 0.000 51.528 0.304 ;
      RECT 51.376 0.000 51.224 0.304 ;
      RECT 51.072 0.000 50.920 0.304 ;
      RECT 49.856 0.000 49.704 0.304 ;
      RECT 48.640 0.000 48.488 0.304 ;
      RECT 47.424 0.000 47.272 0.304 ;
      RECT 46.208 0.000 46.056 0.304 ;
      RECT 44.992 0.000 44.840 0.304 ;
      RECT 43.776 0.000 43.624 0.304 ;
      RECT 42.560 0.000 42.408 0.304 ;
      RECT 41.344 0.000 41.192 0.304 ;
      RECT 40.128 0.000 39.976 0.304 ;
      RECT 38.912 0.000 38.760 0.304 ;
      RECT 37.696 0.000 37.544 0.304 ;
      RECT 36.480 0.000 36.328 0.304 ;
      RECT 35.264 0.000 35.112 0.304 ;
      RECT 34.048 0.000 33.896 0.304 ;
      RECT 32.832 0.000 32.680 0.304 ;
      RECT 54.960 46.056 55.264 50.136 ;
      RECT 54.960 42.408 55.264 45.600 ;
      RECT 54.960 38.760 55.264 41.952 ;
      RECT 54.960 35.112 55.264 38.304 ;
      RECT 54.960 31.464 55.264 34.656 ;
      RECT 54.960 13.376 55.264 31.008 ;
      RECT 54.960 0.304 55.264 12.920 ;
      RECT 0.000 0.000 3.432 0.304 ;
      RECT 3.888 0.000 3.736 0.304 ;
      RECT 4.192 0.000 4.040 0.304 ;
      RECT 5.408 0.000 5.256 0.304 ;
      RECT 6.624 0.000 6.472 0.304 ;
      RECT 7.840 0.000 7.688 0.304 ;
      RECT 9.056 0.000 8.904 0.304 ;
      RECT 10.272 0.000 10.120 0.304 ;
      RECT 11.488 0.000 11.336 0.304 ;
      RECT 12.704 0.000 12.552 0.304 ;
      RECT 13.920 0.000 13.768 0.304 ;
      RECT 15.136 0.000 14.984 0.304 ;
      RECT 16.352 0.000 16.200 0.304 ;
      RECT 17.568 0.000 17.416 0.304 ;
      RECT 18.784 0.000 18.632 0.304 ;
      RECT 20.000 0.000 19.848 0.304 ;
      RECT 21.216 0.000 21.064 0.304 ;
      RECT 22.432 0.000 22.280 0.304 ;
      RECT 23.648 0.000 31.464 0.304 ;
      RECT 0.000 46.056 0.304 50.136 ;
      RECT 0.000 42.408 0.304 45.600 ;
      RECT 0.000 38.760 0.304 41.952 ;
      RECT 0.000 35.112 0.304 38.304 ;
      RECT 0.000 31.464 0.304 34.656 ;
      RECT 0.000 13.376 0.304 31.008 ;
      RECT 0.000 0.304 0.304 12.920 ;
      RECT 0.000 50.136 5.043 52.288 ;
      RECT 7.355 50.136 7.763 52.288 ;
      RECT 10.067 50.136 55.264 52.288 ;
      RECT 0.304 0.304 54.960 50.136 ;
  END

END sram8t17x64

END LIBRARY
